module radixSort(inArray);
  input [1023:0] inArray;

endmodule

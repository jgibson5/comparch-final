module radixSort()

endmodule

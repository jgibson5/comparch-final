module bubble (inArray);
{
    
  
  
}

